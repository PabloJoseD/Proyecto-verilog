/*  Circuitos Digitales 1
    I ciclo 2022  
Autor: Pablo Duran Segura */

//El presente programa describe un módulo COMPARATOR que compara las magnitudes de 2 bits por medio de dos multiplexores 

`include "MUX4x1_Case.v"    //se incluye el archivo del MUX4x1 para luego instanciarlo

module  COMPARATOR( input A,B,   //entradas, cada una de 1 bit
                 output K,L);  //salidas, cada una de 1 bit

reg [3:0]  I;

//instancio el modulo MUX para definir las entradas, lineas de seleccion y salidas diseñadas con los mapas de Karnaugh y las tablas de verdad
MUX4x1_Case MuxK (.I({1,0,1,1}), .S({A,B}), Y.(K)); //multiplexor que resuelve K
MUX4x1_Case MuxL (.I({1,1,0,1}), .S({A,B}), Y.(K));  //multiplexor que resuelve L
  

endmodule   
